* Extracted by KLayout with SG13G2 LVS runset on : 28/01/2026 01:08

.SUBCKT DLINE VSS A Y VIN VDD|VOUT
M$1 \$2 VIN VSS VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p AD=0.1428p PS=1.52u
+ PD=1.1u
M$2 VSS \$2 \$3 VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p AD=0.1428p PS=1.1u
+ PD=1.52u
M$3 \$5 VIN VSS VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p AD=0.1428p PS=1.52u
+ PD=1.1u
M$4 VSS \$5 \$6 VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p AD=0.1428p PS=1.1u
+ PD=1.52u
M$5 VSS \$3 \$11 VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1405p AD=0.2373p
+ PS=1.15u PD=1.97u
M$6 VSS \$11 \$4 VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1405p AD=0.2516p
+ PS=1.15u PD=2.16u
M$7 VSS \$6 \$12 VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1405p AD=0.2373p
+ PS=1.15u PD=1.97u
M$8 VSS \$12 \$4 VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1405p AD=0.2516p
+ PS=1.15u PD=2.16u
M$9 VSS \$4 \$7 VSS sg13_lv_nmos L=0.13u W=2.96u AS=0.6734p AD=0.6734p PS=5.52u
+ PD=5.52u
M$13 VSS \$7 A VSS sg13_lv_nmos L=0.13u W=5.92u AS=1.2395p AD=1.2395p PS=10.01u
+ PD=10.01u
M$21 VSS A Y VSS sg13_lv_nmos L=0.13u W=11.84u AS=2.3606p AD=2.3606p PS=18.96u
+ PD=18.96u
M$37 VDD|VOUT VIN \$2 VDD|VOUT sg13_lv_pmos L=0.13u W=0.42u AS=0.2931p
+ AD=0.1428p PS=1.65u PD=1.52u
M$38 VDD|VOUT \$2 \$3 VDD|VOUT sg13_lv_pmos L=0.13u W=1u AS=0.2931p AD=0.37p
+ PS=1.65u PD=2.74u
M$39 VDD|VOUT VIN \$5 VDD|VOUT sg13_lv_pmos L=0.13u W=0.42u AS=0.2931p
+ AD=0.1428p PS=1.65u PD=1.52u
M$40 VDD|VOUT \$5 \$6 VDD|VOUT sg13_lv_pmos L=0.13u W=1u AS=0.2931p AD=0.37p
+ PS=1.65u PD=2.74u
M$41 \$11 \$3 VDD|VOUT VDD|VOUT sg13_lv_pmos L=0.13u W=1u AS=0.565p AD=0.2245p
+ PS=3.13u PD=1.53u
M$42 VDD|VOUT \$11 \$4 VDD|VOUT sg13_lv_pmos L=0.13u W=1.12u AS=0.2245p
+ AD=0.3808p PS=1.53u PD=2.92u
M$43 \$12 \$6 VDD|VOUT VDD|VOUT sg13_lv_pmos L=0.13u W=1u AS=0.565p AD=0.2245p
+ PS=3.13u PD=1.53u
M$44 VDD|VOUT \$12 \$4 VDD|VOUT sg13_lv_pmos L=0.13u W=1.12u AS=0.2245p
+ AD=0.3808p PS=1.53u PD=2.92u
M$45 VDD|VOUT \$4 \$7 VDD|VOUT sg13_lv_pmos L=0.13u W=4.48u AS=1.0192p
+ AD=1.0192p PS=7.42u PD=7.42u
M$49 VDD|VOUT \$7 A VDD|VOUT sg13_lv_pmos L=0.13u W=8.96u AS=1.876p AD=1.876p
+ PS=13.43u PD=13.43u
M$57 VDD|VOUT A Y VDD|VOUT sg13_lv_pmos L=0.13u W=17.92u AS=3.6288p AD=3.5728p
+ PS=25.52u PD=25.42u
.ENDS DLINE
